library verilog;
use verilog.vl_types.all;
entity a25_decode is
    port(
        quick_n_reset   : in     vl_logic;
        i_clk           : in     vl_logic;
        i_fetch_instruction: in     vl_logic_vector(31 downto 0);
        i_access_stall  : in     vl_logic;
        i_irq           : in     vl_logic;
        i_firq          : in     vl_logic;
        i_dabt          : in     vl_logic;
        i_iabt          : in     vl_logic;
        i_adex          : in     vl_logic;
        i_execute_iaddress: in     vl_logic_vector(31 downto 0);
        i_execute_daddress: in     vl_logic_vector(31 downto 0);
        i_abt_status    : in     vl_logic_vector(7 downto 0);
        i_execute_status_bits: in     vl_logic_vector(31 downto 0);
        i_multiply_done : in     vl_logic;
        o_imm32         : out    vl_logic_vector(31 downto 0);
        o_imm_shift_amount: out    vl_logic_vector(4 downto 0);
        o_shift_imm_zero: out    vl_logic;
        o_condition     : out    vl_logic_vector(3 downto 0);
        o_decode_exclusive: out    vl_logic;
        o_decode_iaccess: out    vl_logic;
        o_decode_daccess: out    vl_logic;
        o_status_bits_mode: out    vl_logic_vector(1 downto 0);
        o_status_bits_irq_mask: out    vl_logic;
        o_status_bits_firq_mask: out    vl_logic;
        o_rm_sel        : out    vl_logic_vector(3 downto 0);
        o_rs_sel        : out    vl_logic_vector(3 downto 0);
        o_load_rd       : out    vl_logic_vector(7 downto 0);
        o_rn_sel        : out    vl_logic_vector(3 downto 0);
        o_barrel_shift_amount_sel: out    vl_logic_vector(1 downto 0);
        o_barrel_shift_data_sel: out    vl_logic_vector(1 downto 0);
        o_barrel_shift_function: out    vl_logic_vector(1 downto 0);
        o_alu_function  : out    vl_logic_vector(8 downto 0);
        o_multiply_function: out    vl_logic_vector(1 downto 0);
        o_interrupt_vector_sel: out    vl_logic_vector(2 downto 0);
        o_iaddress_sel  : out    vl_logic_vector(3 downto 0);
        o_daddress_sel  : out    vl_logic_vector(3 downto 0);
        o_pc_sel        : out    vl_logic_vector(2 downto 0);
        o_byte_enable_sel: out    vl_logic_vector(1 downto 0);
        o_status_bits_sel: out    vl_logic_vector(2 downto 0);
        o_reg_write_sel : out    vl_logic_vector(2 downto 0);
        o_user_mode_regs_store_nxt: out    vl_logic;
        o_firq_not_user_mode: out    vl_logic;
        o_write_data_wen: out    vl_logic;
        o_base_address_wen: out    vl_logic;
        o_pc_wen        : out    vl_logic;
        o_reg_bank_wen  : out    vl_logic_vector(14 downto 0);
        o_status_bits_flags_wen: out    vl_logic;
        o_status_bits_mode_wen: out    vl_logic;
        o_status_bits_irq_mask_wen: out    vl_logic;
        o_status_bits_firq_mask_wen: out    vl_logic;
        o_copro_opcode1 : out    vl_logic_vector(2 downto 0);
        o_copro_opcode2 : out    vl_logic_vector(2 downto 0);
        o_copro_crn     : out    vl_logic_vector(3 downto 0);
        o_copro_crm     : out    vl_logic_vector(3 downto 0);
        o_copro_num     : out    vl_logic_vector(3 downto 0);
        o_copro_operation: out    vl_logic_vector(1 downto 0);
        o_copro_write_data_wen: out    vl_logic;
        o_iabt_trigger  : out    vl_logic;
        o_iabt_address  : out    vl_logic_vector(31 downto 0);
        o_iabt_status   : out    vl_logic_vector(7 downto 0);
        o_dabt_trigger  : out    vl_logic;
        o_dabt_address  : out    vl_logic_vector(31 downto 0);
        o_dabt_status   : out    vl_logic_vector(7 downto 0);
        o_conflict      : out    vl_logic;
        o_rn_use_read   : out    vl_logic;
        o_rm_use_read   : out    vl_logic;
        o_rs_use_read   : out    vl_logic;
        o_rd_use_read   : out    vl_logic
    );
end a25_decode;
