library verilog;
use verilog.vl_types.all;
entity a25_execute is
    port(
        quick_n_reset   : in     vl_logic;
        i_clk           : in     vl_logic;
        i_access_stall  : in     vl_logic;
        i_mem_stall     : in     vl_logic;
        i_wb_read_data  : in     vl_logic_vector(31 downto 0);
        i_wb_read_data_valid: in     vl_logic;
        i_wb_load_rd    : in     vl_logic_vector(9 downto 0);
        i_copro_read_data: in     vl_logic_vector(31 downto 0);
        i_decode_iaccess: in     vl_logic;
        i_decode_daccess: in     vl_logic;
        i_decode_load_rd: in     vl_logic_vector(7 downto 0);
        o_copro_write_data: out    vl_logic_vector(31 downto 0);
        o_write_data    : out    vl_logic_vector(31 downto 0);
        o_iaddress      : out    vl_logic_vector(31 downto 0);
        o_iaddress_nxt  : out    vl_logic_vector(31 downto 0);
        o_iaddress_valid: out    vl_logic;
        o_daddress      : out    vl_logic_vector(31 downto 0);
        o_daddress_nxt  : out    vl_logic_vector(31 downto 0);
        o_daddress_valid: out    vl_logic;
        o_adex          : out    vl_logic;
        o_priviledged   : out    vl_logic;
        o_exclusive     : out    vl_logic;
        o_write_enable  : out    vl_logic;
        o_byte_enable   : out    vl_logic_vector(3 downto 0);
        o_exec_load_rd  : out    vl_logic_vector(7 downto 0);
        o_status_bits   : out    vl_logic_vector(31 downto 0);
        o_multiply_done : out    vl_logic;
        i_status_bits_mode: in     vl_logic_vector(1 downto 0);
        i_status_bits_irq_mask: in     vl_logic;
        i_status_bits_firq_mask: in     vl_logic;
        i_imm32         : in     vl_logic_vector(31 downto 0);
        i_imm_shift_amount: in     vl_logic_vector(4 downto 0);
        i_shift_imm_zero: in     vl_logic;
        i_condition     : in     vl_logic_vector(3 downto 0);
        i_decode_exclusive: in     vl_logic;
        i_rm_sel        : in     vl_logic_vector(3 downto 0);
        i_rs_sel        : in     vl_logic_vector(3 downto 0);
        i_rn_sel        : in     vl_logic_vector(3 downto 0);
        i_barrel_shift_amount_sel: in     vl_logic_vector(1 downto 0);
        i_barrel_shift_data_sel: in     vl_logic_vector(1 downto 0);
        i_barrel_shift_function: in     vl_logic_vector(1 downto 0);
        i_alu_function  : in     vl_logic_vector(8 downto 0);
        i_multiply_function: in     vl_logic_vector(1 downto 0);
        i_interrupt_vector_sel: in     vl_logic_vector(2 downto 0);
        i_iaddress_sel  : in     vl_logic_vector(3 downto 0);
        i_daddress_sel  : in     vl_logic_vector(3 downto 0);
        i_pc_sel        : in     vl_logic_vector(2 downto 0);
        i_byte_enable_sel: in     vl_logic_vector(1 downto 0);
        i_status_bits_sel: in     vl_logic_vector(2 downto 0);
        i_reg_write_sel : in     vl_logic_vector(2 downto 0);
        i_user_mode_regs_store_nxt: in     vl_logic;
        i_firq_not_user_mode: in     vl_logic;
        i_write_data_wen: in     vl_logic;
        i_base_address_wen: in     vl_logic;
        i_pc_wen        : in     vl_logic;
        i_reg_bank_wen  : in     vl_logic_vector(14 downto 0);
        i_status_bits_flags_wen: in     vl_logic;
        i_status_bits_mode_wen: in     vl_logic;
        i_status_bits_irq_mask_wen: in     vl_logic;
        i_status_bits_firq_mask_wen: in     vl_logic;
        i_copro_write_data_wen: in     vl_logic;
        i_conflict      : in     vl_logic;
        i_rn_use_read   : in     vl_logic;
        i_rm_use_read   : in     vl_logic;
        i_rs_use_read   : in     vl_logic;
        i_rd_use_read   : in     vl_logic;
        status_bits_mode: out    vl_logic_vector(1 downto 0);
        status_bits_flags: out    vl_logic_vector(3 downto 0);
        status_bits_irq_mask: out    vl_logic;
        status_bits_firq_mask: out    vl_logic
    );
end a25_execute;
