library verilog;
use verilog.vl_types.all;
entity dumpvcd is
end dumpvcd;
