library verilog;
use verilog.vl_types.all;
entity a25_register_bank is
    port(
        quick_n_reset   : in     vl_logic;
        i_clk           : in     vl_logic;
        i_access_stall  : in     vl_logic;
        i_mem_stall     : in     vl_logic;
        i_mode_idec     : in     vl_logic_vector(1 downto 0);
        i_mode_exec     : in     vl_logic_vector(1 downto 0);
        i_mode_rds_exec : in     vl_logic_vector(3 downto 0);
        i_firq_not_user_mode: in     vl_logic;
        i_rm_sel        : in     vl_logic_vector(3 downto 0);
        i_rs_sel        : in     vl_logic_vector(3 downto 0);
        i_rn_sel        : in     vl_logic_vector(3 downto 0);
        i_pc_wen        : in     vl_logic;
        i_reg_bank_wen  : in     vl_logic_vector(14 downto 0);
        i_pc            : in     vl_logic_vector(23 downto 0);
        i_reg           : in     vl_logic_vector(31 downto 0);
        i_wb_read_data  : in     vl_logic_vector(31 downto 0);
        i_wb_read_data_valid: in     vl_logic;
        i_wb_read_data_rd: in     vl_logic_vector(3 downto 0);
        i_wb_user_mode  : in     vl_logic;
        i_status_bits_flags: in     vl_logic_vector(3 downto 0);
        i_status_bits_irq_mask: in     vl_logic;
        i_status_bits_firq_mask: in     vl_logic;
        o_rm            : out    vl_logic_vector(31 downto 0);
        o_rs            : out    vl_logic_vector(31 downto 0);
        o_rd            : out    vl_logic_vector(31 downto 0);
        o_rn            : out    vl_logic_vector(31 downto 0);
        o_pc            : out    vl_logic_vector(31 downto 0);
        r0_out          : out    vl_logic_vector(31 downto 0);
        r1_out          : out    vl_logic_vector(31 downto 0);
        r2_out          : out    vl_logic_vector(31 downto 0);
        r3_out          : out    vl_logic_vector(31 downto 0);
        r4_out          : out    vl_logic_vector(31 downto 0);
        r5_out          : out    vl_logic_vector(31 downto 0);
        r6_out          : out    vl_logic_vector(31 downto 0);
        r7_out          : out    vl_logic_vector(31 downto 0);
        r8_out          : out    vl_logic_vector(31 downto 0);
        r9_out          : out    vl_logic_vector(31 downto 0);
        r10_out         : out    vl_logic_vector(31 downto 0);
        r11_out         : out    vl_logic_vector(31 downto 0);
        r12_out         : out    vl_logic_vector(31 downto 0);
        r13_out         : out    vl_logic_vector(31 downto 0);
        r14_out         : out    vl_logic_vector(31 downto 0);
        r15_out_rm      : out    vl_logic_vector(31 downto 0);
        r15_out_rn      : out    vl_logic_vector(31 downto 0);
        r14_svc         : out    vl_logic_vector(31 downto 0);
        r14_irq         : out    vl_logic_vector(31 downto 0);
        r14_firq        : out    vl_logic_vector(31 downto 0);
        r0              : out    vl_logic_vector(31 downto 0);
        r1              : out    vl_logic_vector(31 downto 0);
        r2              : out    vl_logic_vector(31 downto 0);
        r3              : out    vl_logic_vector(31 downto 0);
        r4              : out    vl_logic_vector(31 downto 0);
        r5              : out    vl_logic_vector(31 downto 0);
        r6              : out    vl_logic_vector(31 downto 0);
        r7              : out    vl_logic_vector(31 downto 0);
        r8              : out    vl_logic_vector(31 downto 0);
        r9              : out    vl_logic_vector(31 downto 0);
        r10             : out    vl_logic_vector(31 downto 0);
        r11             : out    vl_logic_vector(31 downto 0);
        r12             : out    vl_logic_vector(31 downto 0);
        r13             : out    vl_logic_vector(31 downto 0);
        r14             : out    vl_logic_vector(31 downto 0);
        r15             : out    vl_logic_vector(23 downto 0)
    );
end a25_register_bank;
